module GoldenSnitch(
    clk,
    rst,
    im_addr,
    im_DI,
    dm_web,
    dm_addr,
    dm_DI,
    dm_DO
);








endmodule

