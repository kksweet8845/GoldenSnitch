module MainCtrl(
    opcode,
    funct3,
    funct7,

);







endmodule