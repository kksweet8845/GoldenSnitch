module GS_Core
    import gs_pkg::*
#(
    BOOT_ADDR       = 0,
    ADDR_SIZE       = 32,
    WORD_SIZE       = 32,
    BYTES           = 4 
)
(
    input   logic           clk,
    input   logic           rst,
    //* Instr memory
    output  logic   [ADDR_SIZE-1:0] im_addr_o,
    input   logic   [WORD_SIZE-1:0] im_data_i,

    //* Data memory
    output  logic   [ADDR_SIZE-1:0] dm_addr_o,
    input   logic   [WORD_SIZE-1:0] dm_data_i,
    output  logic   [WORD_SIZE-1:0] dm_data_o,
    output  logic   [BYTES-1:0]     dm_web
);


/*=============================================================================+
/        // ██╗███████╗    ░██████╗████████╗░█████╗░░██████╗░███████╗        /
/        // ██║██╔════╝    ██╔════╝╚══██╔══╝██╔══██╗██╔════╝░██╔════╝        /
/        // ██║█████╗░░    ╚█████╗░░░░██║░░░███████║██║░░██╗░█████╗░░        /
/        // ██║██╔══╝░░    ░╚═══██╗░░░██║░░░██╔══██║██║░░╚██╗██╔══╝░░        /
/        // ██║██║░░░░░    ██████╔╝░░░██║░░░██║░░██║╚██████╔╝███████╗        /
/        // ╚═╝╚═╝░░░░░    ╚═════╝░░░░╚═╝░░░╚═╝░░╚═╝░╚═════╝░╚══════╝        /
 +=============================================================================*/













/*=============================================================================+
/          ██╗██████╗░    ░██████╗████████╗░█████╗░░██████╗░███████╗           /
/          ██║██╔══██╗    ██╔════╝╚══██╔══╝██╔══██╗██╔════╝░██╔════╝           /
/          ██║██║░░██║    ╚█████╗░░░░██║░░░███████║██║░░██╗░█████╗░░           /
/          ██║██║░░██║    ░╚═══██╗░░░██║░░░██╔══██║██║░░╚██╗██╔══╝░░           /
/          ██║██████╔╝    ██████╔╝░░░██║░░░██║░░██║╚██████╔╝███████╗           /
/          ╚═╝╚═════╝░    ╚═════╝░░░░╚═╝░░░╚═╝░░╚═╝░╚═════╝░╚══════╝           /
 +=============================================================================*/



/*=============================================================================+
/        ███████╗██╗░░██╗    ░██████╗████████╗░█████╗░░██████╗░███████╗        /
/        ██╔════╝╚██╗██╔╝    ██╔════╝╚══██╔══╝██╔══██╗██╔════╝░██╔════╝        /
/        █████╗░░░╚███╔╝░    ╚█████╗░░░░██║░░░███████║██║░░██╗░█████╗░░        /
/        ██╔══╝░░░██╔██╗░    ░╚═══██╗░░░██║░░░██╔══██║██║░░╚██╗██╔══╝░░        /
/        ███████╗██╔╝╚██╗    ██████╔╝░░░██║░░░██║░░██║╚██████╔╝███████╗        /
/        ╚══════╝╚═╝░░╚═╝    ╚═════╝░░░░╚═╝░░░╚═╝░░╚═╝░╚═════╝░╚══════╝        /
 +=============================================================================*/





/*=============================================================================+
/     ░██╗░░░░░░░██╗██████╗░    ░██████╗████████╗░█████╗░░██████╗░███████╗     /
/     ░██║░░██╗░░██║██╔══██╗    ██╔════╝╚══██╔══╝██╔══██╗██╔════╝░██╔════╝     /
/     ░╚██╗████╗██╔╝██████╦╝    ╚█████╗░░░░██║░░░███████║██║░░██╗░█████╗░░     /
/     ░░████╔═████║░██╔══██╗    ░╚═══██╗░░░██║░░░██╔══██║██║░░╚██╗██╔══╝░░     /
/     ░░╚██╔╝░╚██╔╝░██████╦╝    ██████╔╝░░░██║░░░██║░░██║╚██████╔╝███████╗     /
/     ░░░╚═╝░░░╚═╝░░╚═════╝░    ╚═════╝░░░░╚═╝░░░╚═╝░░╚═╝░╚═════╝░╚══════╝     /
 +=============================================================================*/
















































endmodule